VERSION 5.8 ;

MACRO analog_blockage
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN analog_blockage 0 0 ;
  SIZE 584.0 BY 260.0 ;

  OBS
    LAYER TopMetal2 ;
      RECT 0 0 584.0 260.0 ;
  END
  OBS
    LAYER TopMetal1 ;
      RECT 0 0 584.0 260.0 ;
  END
  OBS
    LAYER Metal5 ;
      RECT 0 0 584.0 260.0 ;
  END
END analog_blockage